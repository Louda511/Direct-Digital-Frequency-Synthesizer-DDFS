library ieee;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;



entity LUT_DDFS is
	port (
		LUT_line : in  std_logic_vector(7 downto 0);
		LUT_data : out std_logic_vector(7 downto 0) 
	);
end LUT_DDFS;

architecture rtl of LUT_DDFS is
	type LUT_t is array (natural range 0 to 255) of integer;
	constant LUT: LUT_t := (
		0 => 127,
		1 => 130,
		2 => 133,
		3 => 136,
		4 => 139,
		5 => 142,
		6 => 145,
		7 => 148,
		8 => 151,
		9 => 154,
		10 => 157,
		11 => 160,
		12 => 163,
		13 => 166,
		14 => 169,
		15 => 172,
		16 => 175,
		17 => 178,
		18 => 181,
		19 => 184,
		20 => 186,
		21 => 189,
		22 => 192,
		23 => 194,
		24 => 197,
		25 => 200,
		26 => 202,
		27 => 205,
		28 => 207,
		29 => 209,
		30 => 212,
		31 => 214,
		32 => 216,
		33 => 218,
		34 => 221,
		35 => 223,
		36 => 225,
		37 => 227,
		38 => 229,
		39 => 230,
		40 => 232,
		41 => 234,
		42 => 235,
		43 => 237,
		44 => 239,
		45 => 240,
		46 => 241,
		47 => 243,
		48 => 244,
		49 => 245,
		50 => 246,
		51 => 247,
		52 => 248,
		53 => 249,
		54 => 250,
		55 => 250,
		56 => 251,
		57 => 252,
		58 => 252,
		59 => 253,
		60 => 253,
		61 => 253,
		62 => 253,
		63 => 253,
		64 => 254,
		65 => 253,
		66 => 253,
		67 => 253,
		68 => 253,
		69 => 253,
		70 => 252,
		71 => 252,
		72 => 251,
		73 => 250,
		74 => 250,
		75 => 249,
		76 => 248,
		77 => 247,
		78 => 246,
		79 => 245,
		80 => 244,
		81 => 243,
		82 => 241,
		83 => 240,
		84 => 239,
		85 => 237,
		86 => 235,
		87 => 234,
		88 => 232,
		89 => 230,
		90 => 229,
		91 => 227,
		92 => 225,
		93 => 223,
		94 => 221,
		95 => 218,
		96 => 216,
		97 => 214,
		98 => 212,
		99 => 209,
		100 => 207,
		101 => 205,
		102 => 202,
		103 => 200,
		104 => 197,
		105 => 194,
		106 => 192,
		107 => 189,
		108 => 186,
		109 => 184,
		110 => 181,
		111 => 178,
		112 => 175,
		113 => 172,
		114 => 169,
		115 => 166,
		116 => 163,
		117 => 160,
		118 => 157,
		119 => 154,
		120 => 151,
		121 => 148,
		122 => 145,
		123 => 142,
		124 => 139,
		125 => 136,
		126 => 133,
		127 => 130,
		128 => 127,
		129 => 123,
		130 => 120,
		131 => 117,
		132 => 114,
		133 => 111,
		134 => 108,
		135 => 105,
		136 => 102,
		137 => 99,
		138 => 96,
		139 => 93,
		140 => 90,
		141 => 87,
		142 => 84,
		143 => 81,
		144 => 78,
		145 => 75,
		146 => 72,
		147 => 69,
		148 => 67,
		149 => 64,
		150 => 61,
		151 => 59,
		152 => 56,
		153 => 53,
		154 => 51,
		155 => 48,
		156 => 46,
		157 => 44,
		158 => 41,
		159 => 39,
		160 => 37,
		161 => 35,
		162 => 32,
		163 => 30,
		164 => 28,
		165 => 26,
		166 => 24,
		167 => 23,
		168 => 21,
		169 => 19,
		170 => 18,
		171 => 16,
		172 => 14,
		173 => 13,
		174 => 12,
		175 => 10,
		176 => 9,
		177 => 8,
		178 => 7,
		179 => 6,
		180 => 5,
		181 => 4,
		182 => 3,
		183 => 3,
		184 => 2,
		185 => 1,
		186 => 1,
		187 => 0,
		188 => 0,
		189 => 0,
		190 => 0,
		191 => 0,
		192 => 0,
		193 => 0,
		194 => 0,
		195 => 0,
		196 => 0,
		197 => 0,
		198 => 1,
		199 => 1,
		200 => 2,
		201 => 3,
		202 => 3,
		203 => 4,
		204 => 5,
		205 => 6,
		206 => 7,
		207 => 8,
		208 => 9,
		209 => 10,
		210 => 12,
		211 => 13,
		212 => 14,
		213 => 16,
		214 => 18,
		215 => 19,
		216 => 21,
		217 => 23,
		218 => 24,
		219 => 26,
		220 => 28,
		221 => 30,
		222 => 32,
		223 => 35,
		224 => 37,
		225 => 39,
		226 => 41,
		227 => 44,
		228 => 46,
		229 => 48,
		230 => 51,
		231 => 53,
		232 => 56,
		233 => 59,
		234 => 61,
		235 => 64,
		236 => 67,
		237 => 69,
		238 => 72,
		239 => 75,
		240 => 78,
		241 => 81,
		242 => 84,
		243 => 87,
		244 => 90,
		245 => 93,
		246 => 96,
		247 => 99,
		248 => 102,
		249 => 105,
		250 => 108,
		251 => 111,
		252 => 114,
		253 => 117,
		254 => 120,
		255 => 123
);

begin
	LUT_data <= std_logic_vector(TO_UNSIGNED(LUT(TO_INTEGER(unsigned(LUT_line))), 8));
end rtl;
